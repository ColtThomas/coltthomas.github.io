library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity counter_3to12 is
	
end counter_3to12;

architecture Behavioral of counter_3to12 is

begin


end Behavioral;

